
// This is the start of our actual project. 
module fpga_top();

endmodule 